module mmu(
);

endmodule
